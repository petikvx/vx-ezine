� �  �                                                                                                                                                                                                                                                                                                                                                              B	artles A	nd J	aymes                                                                   P
resent:                                                                                                                                                  Computer Virus Cooler                                                                                                                                                                                                                       �����������������    ��x�x�x�� �                                                     ��  ��   �  �� ��    �x�x�x�x�x x                                                     ��  ����� �� � ��   �=x=x=x�x�x�x                                                     �� �� � � �� � ��   ����y�z�x�x�x                                                     ��  � � � � �  ��   ��x�x�x�x�x�                                                     �����������������   � w w����                                                      ��           ��    ��   ��                                                                                                                                 W
a
t
c
h
 
y
o
u
r
 
c
o
m
p
u
t
e
r
 
g
o
 
u
p
 
i
n
 
b
u
b
b
l
e
s
!
                                                                                                                  T	h	i	s	 	i	s	 	B	a	r	t	l	e	s	 	a	n	d	 	J	a	y	m	e	s	,	 	a	n	d	 	t	h	a	n	k	 	y	o	u	 	f	o	r	 	y	o	u	r	 	s	u	p	p	o	r	t	.	                                                                                                                                                                                                                                                                                                                                         � �  �